-- Implements a simple Nios II system for the DE-series board.
-- Inputs: SW7-0 are parallel port inputs to the Nios II system.
-- CLOCK_50 is the system clock.
-- KEY0 is the active-low system reset.
-- Outputs: LED7-0 are parallel port outputs from the Nios II system.
-- SDRAM ports correspond to the SDRAM signals on the DE-series board.
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;

ENTITY ROBOT IS
PORT (
	SW : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	KEY : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
	CLOCK_50 : IN STD_LOGIC;
	LED : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	DRAM_CLK, DRAM_CKE : OUT STD_LOGIC;
	DRAM_ADDR : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	DRAM_BA : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N, DRAM_WE_N : OUT STD_LOGIC;
	DRAM_DQ : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	DRAM_DQM : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	-- Motor Driver DRV8848 interface
	MTRR_P, MTRR_N : OUT STD_LOGIC;
	MTRL_P, MTRL_N : OUT STD_LOGIC;
	MTR_Sleep_n : OUT STD_LOGIC;
	MTR_Fault_n : IN STD_LOGIC;
	-- Sensor power control (A-Cute Car)
	VCC3P3_PWRON_n : OUT STD_LOGIC;
	IR_LED_ON : OUT STD_LOGIC;
	-- ADC LTC2308 interface
	LTC_ADC_CONVST : OUT STD_LOGIC;
	LTC_ADC_SCK : OUT STD_LOGIC;
	LTC_ADC_SDI : OUT STD_LOGIC;
	LTC_ADC_SDO : IN STD_LOGIC );
END ROBOT;

ARCHITECTURE Structure OF ROBOT IS

COMPONENT nios_system_sdram
PORT (
	clk_clk : IN STD_LOGIC;
	reset_reset_n : IN STD_LOGIC;
	sdram_clk_clk : OUT STD_LOGIC;
	leds_export : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	switches_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	sdram_wire_addr : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	sdram_wire_ba : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	sdram_wire_cas_n : OUT STD_LOGIC;
	sdram_wire_cke : OUT STD_LOGIC;
	sdram_wire_cs_n : OUT STD_LOGIC;
	sdram_wire_dq : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	sdram_wire_dqm : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	sdram_wire_ras_n : OUT STD_LOGIC;
	sdram_wire_we_n : OUT STD_LOGIC;
	motor_right_export : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
	motor_left_export : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
	-- Ground sensors PIOs
	sensor_control_export : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	sensor_status_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	sensor_data0_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	sensor_data1_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	sensor_data2_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	sensor_data3_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	sensor_data4_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	sensor_data5_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	sensor_data6_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0) );
END COMPONENT;

COMPONENT capteurs_sol
PORT (
	clk : IN STD_LOGIC;
	reset_n : IN STD_LOGIC;
	data_capture : IN STD_LOGIC;
	data_readyr : OUT STD_LOGIC;
	data0r : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	data1r : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	data2r : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	data3r : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	data4r : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	data5r : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	data6r : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	ADC_CONVSTr : OUT STD_LOGIC;
	ADC_SCK : OUT STD_LOGIC;
	ADC_SDIr : OUT STD_LOGIC;
	ADC_SDO : IN STD_LOGIC );
END COMPONENT;

COMPONENT PWM_generation
PORT (
	clk, reset_n : IN STD_LOGIC;
	s_writedataR, s_writedataL : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
	dc_motor_p_R, dc_motor_n_R : OUT STD_LOGIC;
	dc_motor_p_L, dc_motor_n_L : OUT STD_LOGIC );
END COMPONENT;

-- Fault signal (not used in this version, just monitored)
signal motor_fault : STD_LOGIC;

-- Internal signals for motor control
signal motor_right_data : STD_LOGIC_VECTOR(13 DOWNTO 0);
signal motor_left_data : STD_LOGIC_VECTOR(13 DOWNTO 0);

-- Internal signals for ground sensors
signal sensor_control_sig : STD_LOGIC_VECTOR(7 DOWNTO 0);
signal sensor_status_sig : STD_LOGIC_VECTOR(7 DOWNTO 0);
signal data_capture_sig : STD_LOGIC;
signal data_ready_sig : STD_LOGIC;
signal data0_sig : STD_LOGIC_VECTOR(7 DOWNTO 0);
signal data1_sig : STD_LOGIC_VECTOR(7 DOWNTO 0);
signal data2_sig : STD_LOGIC_VECTOR(7 DOWNTO 0);
signal data3_sig : STD_LOGIC_VECTOR(7 DOWNTO 0);
signal data4_sig : STD_LOGIC_VECTOR(7 DOWNTO 0);
signal data5_sig : STD_LOGIC_VECTOR(7 DOWNTO 0);
signal data6_sig : STD_LOGIC_VECTOR(7 DOWNTO 0);

-- Clock divider for 2 KHz data_capture signal
-- 50 MHz / 2 KHz = 25000
signal clk_div_counter : INTEGER range 0 to 24999 := 0;
signal data_capture_2khz : STD_LOGIC := '0';

-- Instantiate the Nios II system entity generated by the Qsys tool.
BEGIN
NiosII: nios_system_sdram
PORT MAP (
	clk_clk => CLOCK_50,
	reset_reset_n => KEY(0),
	sdram_clk_clk => DRAM_CLK,
	leds_export => LED,
	switches_export => SW,
	sdram_wire_addr => DRAM_ADDR,
	sdram_wire_ba => DRAM_BA,
	sdram_wire_cas_n => DRAM_CAS_N,
	sdram_wire_cke => DRAM_CKE,
	sdram_wire_cs_n => DRAM_CS_N,
	sdram_wire_dq => DRAM_DQ,
	sdram_wire_dqm => DRAM_DQM,
	sdram_wire_ras_n => DRAM_RAS_N,
	sdram_wire_we_n => DRAM_WE_N,
	motor_right_export => motor_right_data,
	motor_left_export => motor_left_data,
	-- Ground sensors
	sensor_control_export => sensor_control_sig,
	sensor_status_export => sensor_status_sig,
	sensor_data0_export => data0_sig,
	sensor_data1_export => data1_sig,
	sensor_data2_export => data2_sig,
	sensor_data3_export => data3_sig,
	sensor_data4_export => data4_sig,
	sensor_data5_export => data5_sig,
	sensor_data6_export => data6_sig );

-- Extract control and status signals
sensor_status_sig <= "0000000" & data_ready_sig;

-- Generate 2 KHz pulse for data_capture
process(CLOCK_50, KEY(0))
begin
	if KEY(0) = '0' then
		clk_div_counter <= 0;
		data_capture_2khz <= '0';
	elsif rising_edge(CLOCK_50) then
		if clk_div_counter = 24999 then
			clk_div_counter <= 0;
			data_capture_2khz <= NOT data_capture_2khz; -- Toggle at 2 KHz
		else
			clk_div_counter <= clk_div_counter + 1;
		end if;
	end if;
end process;

-- Use 2 KHz signal for data capture
data_capture_sig <= data_capture_2khz;

Capteurs: capteurs_sol
PORT MAP (
	clk => CLOCK_50,
	reset_n => KEY(0),
	data_capture => data_capture_sig,
	data_readyr => data_ready_sig,
	data0r => data0_sig,
	data1r => data1_sig,
	data2r => data2_sig,
	data3r => data3_sig,
	data4r => data4_sig,
	data5r => data5_sig,
	data6r => data6_sig,
	ADC_CONVSTr => LTC_ADC_CONVST,
	ADC_SCK => LTC_ADC_SCK,
	ADC_SDIr => LTC_ADC_SDI,
	ADC_SDO => LTC_ADC_SDO );


-- Instantiate PWM generation for motor control
PWM_Motors: PWM_generation
PORT MAP (
	clk => CLOCK_50,
	reset_n => KEY(0),
	s_writedataR => motor_right_data,
	s_writedataL => motor_left_data,
	dc_motor_p_R => MTRR_P,
	dc_motor_n_R => MTRR_N,
	dc_motor_p_L => MTRL_P,
	dc_motor_n_L => MTRL_N );

-- Motor driver control signals
MTR_Sleep_n <= '1'; -- Enable motor driver (active high)
motor_fault <= MTR_Fault_n; -- Monitor fault signal

-- Sensor power control (A-Cute Car)
VCC3P3_PWRON_n <= '0'; -- Enable 3.3V power for sensors (active low)
IR_LED_ON <= '1'; -- Enable IR LEDs for line sensors

END Structure;