-- Implements a simple Nios II system for the DE-series board.
-- Inputs: SW7-0 are parallel port inputs to the Nios II system.
-- CLOCK_50 is the system clock.
-- KEY0 is the active-low system reset.
-- Outputs: LED7-0 are parallel port outputs from the Nios II system.
-- SDRAM ports correspond to the SDRAM signals on the DE-series board.
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;

ENTITY ROBOT IS
PORT (
	SW : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	KEY : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
	CLOCK_50 : IN STD_LOGIC;
	LED : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	DRAM_CLK, DRAM_CKE : OUT STD_LOGIC;
	DRAM_ADDR : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	DRAM_BA : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N, DRAM_WE_N : OUT STD_LOGIC;
	DRAM_DQ : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	DRAM_DQM : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	-- Motor Driver DRV8848 interface
	MTRR_P, MTRR_N : OUT STD_LOGIC;
	MTRL_P, MTRL_N : OUT STD_LOGIC;
	MTR_Sleep_n : OUT STD_LOGIC;
	MTR_Fault_n : IN STD_LOGIC );
END ROBOT;

ARCHITECTURE Structure OF ROBOT IS

COMPONENT nios_system_sdram
PORT (
	clk_clk : IN STD_LOGIC;
	reset_reset_n : IN STD_LOGIC;
	sdram_clk_clk : OUT STD_LOGIC;
	leds_export : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	switches_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	sdram_wire_addr : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	sdram_wire_ba : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	sdram_wire_cas_n : OUT STD_LOGIC;
	sdram_wire_cke : OUT STD_LOGIC;
	sdram_wire_cs_n : OUT STD_LOGIC;
	sdram_wire_dq : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	sdram_wire_dqm : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	sdram_wire_ras_n : OUT STD_LOGIC;
	sdram_wire_we_n : OUT STD_LOGIC;
	motor_right_export : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
	motor_left_export : OUT STD_LOGIC_VECTOR(13 DOWNTO 0) );
END COMPONENT;


COMPONENT PWM_generation
PORT (
	clk, reset_n : IN STD_LOGIC;
	s_writedataR, s_writedataL : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
	dc_motor_p_R, dc_motor_n_R : OUT STD_LOGIC;
	dc_motor_p_L, dc_motor_n_L : OUT STD_LOGIC );
END COMPONENT;

-- Fault signal (not used in this version, just monitored)
signal motor_fault : STD_LOGIC;

-- Internal signals for motor control
signal motor_right_data : STD_LOGIC_VECTOR(13 DOWNTO 0);
signal motor_left_data : STD_LOGIC_VECTOR(13 DOWNTO 0);

-- Instantiate the Nios II system entity generated by the Qsys tool.
BEGIN
NiosII: nios_system_sdram
PORT MAP (
	clk_clk => CLOCK_50,
	reset_reset_n => KEY(0),
	sdram_clk_clk => DRAM_CLK,
	leds_export => LED,
	switches_export => SW,
	sdram_wire_addr => DRAM_ADDR,
	sdram_wire_ba => DRAM_BA,
	sdram_wire_cas_n => DRAM_CAS_N,
	sdram_wire_cke => DRAM_CKE,
	sdram_wire_cs_n => DRAM_CS_N,
	sdram_wire_dq => DRAM_DQ,
	sdram_wire_dqm => DRAM_DQM,
	sdram_wire_ras_n => DRAM_RAS_N,
	sdram_wire_we_n => DRAM_WE_N,
	motor_right_export => motor_right_data,
	motor_left_export => motor_left_data );

-- Instantiate PWM generation for motor control
PWM_Motors: PWM_generation
PORT MAP (
	clk => CLOCK_50,
	reset_n => KEY(0),
	s_writedataR => motor_right_data,
	s_writedataL => motor_left_data,
	dc_motor_p_R => MTRR_P,
	dc_motor_n_R => MTRR_N,
	dc_motor_p_L => MTRL_P,
	dc_motor_n_L => MTRL_N );

-- Motor driver control signals
MTR_Sleep_n <= '1'; -- Enable motor driver (active high)
motor_fault <= MTR_Fault_n; -- Monitor fault signal

END Structure;
